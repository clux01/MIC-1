`ifndef _mic1_include_
`define _mic1_include_

`define MIC1_PROGRAM "ijvmtest.mem"
`define MIC1_MICROCODE "microcode.mem"
`define CONSTANTPOOL_ADDRESS 'hc3
`define LOCALVARIABLEFRAME_ADDRESS 'hc6
`define STACKPOINTER_ADDRESS 'hd6
`define MEMORY_SIZE 'h106

`endif